entity BCD_Decoder is
	port(ABCD: in bit_vector(3 downto 0);
		F: out bit_vector(6 downto 0));
end BCD_Decoder;

architecture behavioral of BCD_Decoder is
begin
	with (ABCD) select
		F <= "1111110" when "0000",
		 "0110000" when "0001",
		 "1101101" when "0010",
		 "1111001" when "0011",
		 "0110011" when "0100",
		 "1011011" when "0101",
		 "1011111" when "0110",
		 "1110000" when "0111",
		 "1111111" when "1000",
		 "1110011" when "1001",
		 "0000001" when others;
end behavioral;