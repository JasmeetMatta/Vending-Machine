entity test is
--empty
end entity;

architecture bench of test is
component fourPin is 
	port (A: in bit;
		B: in bit;
		C: in bit;
		D: in bit;
		F: out bit);
	end component;
signal a_t, b_t, c_t, d_t, f_t: bit;

begin 

uut: fourPin port map(a_t, b_t, c_t, d_t, f_t);

a_t <= '0', '0' after 20 ns, '0' after 40 ns, '0' after 60 ns, '0' after 80 ns, '0' after 100 ns, '0' after 120 ns, '0' after 140 ns, '1' after 160 ns, '1' after 180 ns, '1' after 200 ns, '1' after 220 ns, '1' after 240 ns, '1' after 260 ns,'1' after 280 ns, '1' after 300 ns;
b_t <= '0', '0' after 20 ns, '0' after 40 ns, '0' after 60 ns, '1' after 80 ns, '1' after 100 ns, '1' after 120 ns, '1' after 140 ns, '0' after 160 ns, '0' after 180 ns, '0' after 200 ns, '0' after 220 ns, '1' after 240 ns, '1' after 260 ns,'1' after 280 ns, '1' after 300 ns;
c_t <= '0', '0' after 20 ns, '1' after 40 ns, '1' after 60 ns, '0' after 80 ns, '0' after 100 ns, '1' after 120 ns, '1' after 140 ns, '0' after 160 ns, '0' after 180 ns, '1' after 200 ns, '1' after 220 ns, '0' after 240 ns, '0' after 260 ns,'1' after 280 ns, '1' after 300 ns;
d_t <= '0', '1' after 20 ns, '0' after 40 ns, '1' after 60 ns, '0' after 80 ns, '1' after 100 ns, '0' after 120 ns, '1' after 140 ns, '0' after 160 ns, '1' after 180 ns, '0' after 200 ns, '1' after 220 ns, '0' after 240 ns, '1' after 260 ns,'0' after 280 ns, '1' after 300 ns;
end;

