-- Jasmeet Singh Matta
-- 2023
-- Hardware Engineering
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

entity Input_Display is
	port ( sw0: in STD_LOGIC_VECTOR(1 downto 0);
		sw1: in STD_LOGIC_VECTOR(3 downto 0);
		ResetBtn: in STD_LOGIC;
		Display: out STD_LOGIC_VECTOR (7 downto 0);
		Clk: in STD_LOGIC;
		An0: out STD_LOGIC_VECTOR ( 7 downto 0));
end Input_Display;

architecture behaviour of Input_Display is
	signal Refresh_counter: STD_LOGIC_VECTOR( 19 downto 0);
	signal Led_activation: STD_LOGIC_VECTOR(2 downto 0);
	signal DataDisp: STD_LOGIC_VECTOR(3 downto 0);
	signal Disp: STD_LOGIC_VECTOR(7 downto 0);
begin
	Refresh: process(Clk ,ResetBtn)
	begin 
   		if(ResetBtn='1') then
        		refresh_counter <= (others => '0');
    		elsif(rising_edge(Clk)) then
        		refresh_counter <= refresh_counter+1;
    		end if;
	end Process;
	Led_activation <= Refresh_counter(19 downto 17);
	DisplayBCD: process(Led_Activation)
	begin 
		Case(Led_activation) is
		when "000" =>
			An0 <= "01111111";
			if(sw0 = "00") then
				DataDisp <= "0000";
			elsif(sw0 = "01") then
				DataDisp <= "1101";
			elsif(sw0 = "10") then
				DataDisp <= "1111";
			elsif(Sw0 = "11") then
				DataDisp <= "1101";
			end if;
		when "001" =>
			An0 <= "10111111";
			if(Sw0 = "11") then
				DataDisp <= "1111";
			end if;
		when"010" =>
			An0 <= "11011111";
			if(sw0 = "01") then
				DataDisp <= "0000";
			elsif(sw0 = "10") then
				DataDisp <= "0000";
			elsif(sw0 = "11") then
				DataDisp <= "0001";
			end if;
		when "011" =>
			An0 <= "11101111";
			if(sw0 = "01") then
				DataDisp <= "0110";
			elsif(sw0 = "10") then
				DataDisp <= "0100";
			elsif(sw0 = "11") then
				DataDisp <= "0000";
			end if;
		when "100" =>
			An0 <= "11110111";
			DataDisp <= "0000"; --change it to Display P
		when "101" =>
			An0 <= "11111101";
			if(sw1 = "0000") then
				DataDisp <= "1010";
			elsif(sw1 = "0001") then
				DataDisp <= "1010";
			elsif(sw1 = "0010") then
				DataDisp <= "1010";
			elsif(sw1 = "0011") then
				DataDisp <= "1010";
			elsif(sw1 = "0100") then
				DataDisp <= "1010";
			elsif(sw1 = "0101") then
				DataDisp <= "1010";
			elsif(sw1 = "0110") then
				DataDisp <= "1011";
			elsif(sw1 = "0111") then
				DataDisp <= "1011";
			elsif(sw1 = "1000") then
				DataDisp <= "1011";
			elsif(sw1 = "1001") then
				DataDisp <= "1011";
			elsif(sw1 = "1010") then
				DataDisp <= "1011";
			elsif(sw1 = "1011") then
				DataDisp <= "1011";
			elsif(sw1 = "1100") then
				DataDisp <= "1011";
			elsif(sw1 = "1101") then
				DataDisp <= "1011";
			elsif(sw1 = "1110") then
				DataDisp <= "1100";
			elsif(sw1 = "1111") then
				DataDisp <= "1100";
			end if;
		when others =>
			An0 <= "11111110";
			if(sw1 = "0000") then
				DataDisp <= "0000";
			elsif(sw1 = "0001") then
				DataDisp <= "0010";
			elsif(sw1 = "0010") then
				DataDisp <= "0100";
			elsif(sw1 = "0011") then
				DataDisp <= "0110";
			elsif(sw1 = "0100") then
				DataDisp <= "0010";
			elsif(sw1 = "0101") then
				DataDisp <= "1000";
			elsif(sw1 = "0110") then
				DataDisp <= "0000";
			elsif(sw1 = "0111") then
				DataDisp <= "0010";
			elsif(sw1 = "1000") then
				DataDisp <= "0000";
			elsif(sw1 = "1001") then
				DataDisp <= "0010";
			elsif(sw1 = "1010") then
				DataDisp <= "0100";
			elsif(sw1 = "1011") then
				DataDisp <= "0110";
			elsif(sw1 = "1100") then
				DataDisp <= "0110";
			elsif(sw1 = "1101") then
				DataDisp <= "1000";
			elsif(sw1 = "1110") then
				DataDisp <= "0000";
			elsif(sw1 = "1111") then
				DataDisp <= "0010";
			end if;
		end case;
	end process;
	CallDisp: process (DataDisp)
	begin
    	case DataDisp is
    		when "0000" => Display <= "00000011"; -- "0"     
    		when "0001" => Display <= "10011111"; -- "1" 
    		when "0010" => Display <= "00100101"; -- "2" 
    		when "0011" => Display <= "00001101"; -- "3" 
    		when "0100" => Display <= "10011001"; -- "4" 
    		when "0101" => Display <= "01001001"; -- "5" 
    		when "0110" => Display <= "01000001"; -- "6" 
    		when "0111" => Display <= "00011111"; -- "7" 
    		when "1000" => Display <= "00000001"; -- "8"     
    		when "1001" => Display <= "00001001"; -- "9" 
    		when "1010" => Display <= "00000010"; -- 0.
    		when "1011" => Display <= "10011110"; -- 1.
    		when "1100" => Display <= "00100100"; -- 2.
    		when "1101" => Display <= "01100011"; -- C
    		when "1110" => Display <= "01100001"; -- E
    		when others => Display <= "01110001"; -- F
    	end case;
	end process;
end;
	
